----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07.10.2019 10:22:29
-- Design Name: 
-- Module Name: sinus_form_generator - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
use IEEE.Numeric_Std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sinus_form_generator is
    Port ( 
      clk   : in std_logic;
      rst   : in std_logic;
      start : in std_logic;
      addr  : out std_logic_vector(10 downto 0);
      data  : out std_logic_vector(7 downto 0);
      wr_en : out std_logic
    );
end sinus_form_generator;

architecture Behavioral of sinus_form_generator is
    type sin_form_ROM   is array (0 to 2047) of std_logic_vector(7 downto 0);
    constant sin_form : sin_form_ROM :=
    (x"7F",
     x"7F",
     x"80",
     x"80",
     x"81",
     x"81",
     x"81",
     x"82",
     x"82",
     x"82",
     x"83",
     x"83",
     x"84",
     x"84",
     x"84",
     x"85",
     x"85",
     x"85",
     x"86",
     x"86",
     x"87",
     x"87",
     x"87",
     x"7E",
     x"88",
     x"88",
     x"89",
     x"89",
     x"89",
     x"8A",
     x"8A",
     x"8A",
     x"8B",
     x"8B",
     x"8C",
     x"8C",
     x"8C",
     x"8D",
     x"8D",
     x"8D",
     x"8E",
     x"8E",
     x"8F",
     x"8F",
     x"8F",
     x"90",
     x"90",
     x"90",
     x"91",
     x"91",
     x"92",
     x"92",
     x"92",
     x"93",
     x"93",
     x"93",
     x"94",
     x"94",
     x"95",
     x"95",
     x"95",
     x"96",
     x"96",
     x"96",
     x"97",
     x"97",
     x"98",
     x"98",
     x"98",
     x"99",
     x"99",
     x"99",
     x"9A",
     x"9A",
     x"9B",
     x"9B",
     x"9B",
     x"9C",
     x"9C",
     x"9C",
     x"9D",
     x"9D",
     x"9D",
     x"9E",
     x"9E",
     x"9F",
     x"9F",
     x"9F",
     x"A0",
     x"A0",
     x"A0",
     x"A1",
     x"A1",
     x"A2",
     x"A2",
     x"A2",
     x"A3",
     x"A3",
     x"A3",
     x"A4",
     x"A4",
     x"A4",
     x"A5",
     x"A5",
     x"A6",
     x"A6",
     x"A6",
     x"A7",
     x"A7",
     x"A7",
     x"A8",
     x"A8",
     x"A8",
     x"A9",
     x"A9",
     x"A9",
     x"AA",
     x"AA",
     x"AB",
     x"AB",
     x"AB",
     x"AC",
     x"AC",
     x"AC",
     x"AD",
     x"AD",
     x"AD",
     x"AE",
     x"AE",
     x"AE",
     x"AF",
     x"AF",
     x"B0",
     x"B0",
     x"B0",
     x"B1",
     x"B1",
     x"B1",
     x"B2",
     x"B2",
     x"B2",
     x"B3",
     x"B3",
     x"B3",
     x"B4",
     x"B4",
     x"B4",
     x"B5",
     x"B5",
     x"B5",
     x"B6",
     x"B6",
     x"B6",
     x"B7",
     x"B7",
     x"B7",
     x"B8",
     x"B8",
     x"B8",
     x"B9",
     x"B9",
     x"B9",
     x"BA",
     x"BA",
     x"BA",
     x"BB",
     x"BB",
     x"BB",
     x"BC",
     x"BC",
     x"BC",
     x"BD",
     x"BD",
     x"BD",
     x"BE",
     x"BE",
     x"BE",
     x"BF",
     x"BF",
     x"BF",
     x"C0",
     x"C0",
     x"C0",
     x"C1",
     x"C1",
     x"C1",
     x"C2",
     x"C2",
     x"C2",
     x"C3",
     x"C3",
     x"C3",
     x"C4",
     x"C4",
     x"C4",
     x"C5",
     x"C5",
     x"C5",
     x"C5",
     x"C6",
     x"C6",
     x"C6",
     x"C7",
     x"C7",
     x"C7",
     x"C8",
     x"C8",
     x"C8",
     x"C9",
     x"C9",
     x"C9",
     x"C9",
     x"CA",
     x"CA",
     x"CA",
     x"CB",
     x"CB",
     x"CB",
     x"CC",
     x"CC",
     x"CC",
     x"CC",
     x"CD",
     x"CD",
     x"CD",
     x"CE",
     x"CE",
     x"CE",
     x"CF",
     x"CF",
     x"CF",
     x"CF",
     x"D0",
     x"D0",
     x"D0",
     x"D1",
     x"D1",
     x"D1",
     x"D1",
     x"D2",
     x"D2",
     x"D2",
     x"D3",
     x"D3",
     x"D3",
     x"D3",
     x"D4",
     x"D4",
     x"D4",
     x"D5",
     x"D5",
     x"D5",
     x"D5",
     x"D6",
     x"D6",
     x"D6",
     x"D6",
     x"D7",
     x"D7",
     x"D7",
     x"D7",
     x"D8",
     x"D8",
     x"D8",
     x"D9",
     x"D9",
     x"D9",
     x"D9",
     x"DA",
     x"DA",
     x"DA",
     x"DA",
     x"DB",
     x"DB",
     x"DB",
     x"DB",
     x"DC",
     x"DC",
     x"DC",
     x"DC",
     x"DD",
     x"DD",
     x"DD",
     x"DD",
     x"DE",
     x"DE",
     x"DE",
     x"DE",
     x"DF",
     x"DF",
     x"DF",
     x"DF",
     x"E0",
     x"E0",
     x"E0",
     x"E0",
     x"E1",
     x"E1",
     x"E1",
     x"E1",
     x"E1",
     x"E2",
     x"E2",
     x"E2",
     x"E2",
     x"E3",
     x"E3",
     x"E3",
     x"E3",
     x"E3",
     x"E4",
     x"E4",
     x"E4",
     x"E4",
     x"E5",
     x"E5",
     x"E5",
     x"E5",
     x"E5",
     x"E6",
     x"E6",
     x"E6",
     x"E6",
     x"E7",
     x"E7",
     x"E7",
     x"E7",
     x"E7",
     x"E8",
     x"E8",
     x"E8",
     x"E8",
     x"E8",
     x"E9",
     x"E9",
     x"E9",
     x"E9",
     x"E9",
     x"EA",
     x"EA",
     x"EA",
     x"EA",
     x"EA",
     x"EB",
     x"EB",
     x"EB",
     x"EB",
     x"EB",
     x"EB",
     x"EC",
     x"EC",
     x"EC",
     x"EC",
     x"EC",
     x"ED",
     x"ED",
     x"ED",
     x"ED",
     x"ED",
     x"ED",
     x"EE",
     x"EE",
     x"EE",
     x"EE",
     x"EE",
     x"EE",
     x"EF",
     x"EF",
     x"EF",
     x"EF",
     x"EF",
     x"EF",
     x"F0",
     x"F0",
     x"F0",
     x"F0",
     x"F0",
     x"F0",
     x"F1",
     x"F1",
     x"F1",
     x"F1",
     x"F1",
     x"F1",
     x"F1",
     x"F2",
     x"F2",
     x"F2",
     x"F2",
     x"F2",
     x"F2",
     x"F2",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F4",
     x"F4",
     x"F4",
     x"F4",
     x"F4",
     x"F4",
     x"F4",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FB",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"FA",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F9",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F8",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F7",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F6",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F5",
     x"F4",
     x"F4",
     x"F4",
     x"F4",
     x"F4",
     x"F4",
     x"F4",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F3",
     x"F2",
     x"F2",
     x"F2",
     x"F2",
     x"F2",
     x"F2",
     x"F2",
     x"F1",
     x"F1",
     x"F1",
     x"F1",
     x"F1",
     x"F1",
     x"F1",
     x"F0",
     x"F0",
     x"F0",
     x"F0",
     x"F0",
     x"F0",
     x"EF",
     x"EF",
     x"EF",
     x"EF",
     x"EF",
     x"EF",
     x"EE",
     x"EE",
     x"EE",
     x"EE",
     x"EE",
     x"EE",
     x"ED",
     x"ED",
     x"ED",
     x"ED",
     x"ED",
     x"ED",
     x"EC",
     x"EC",
     x"EC",
     x"EC",
     x"EC",
     x"EB",
     x"EB",
     x"EB",
     x"EB",
     x"EB",
     x"EB",
     x"EA",
     x"EA",
     x"EA",
     x"EA",
     x"EA",
     x"E9",
     x"E9",
     x"E9",
     x"E9",
     x"E9",
     x"E8",
     x"E8",
     x"E8",
     x"E8",
     x"E8",
     x"E7",
     x"E7",
     x"E7",
     x"E7",
     x"E7",
     x"E6",
     x"E6",
     x"E6",
     x"E6",
     x"E5",
     x"E5",
     x"E5",
     x"E5",
     x"E5",
     x"E4",
     x"E4",
     x"E4",
     x"E4",
     x"E3",
     x"E3",
     x"E3",
     x"E3",
     x"E3",
     x"E2",
     x"E2",
     x"E2",
     x"E2",
     x"E1",
     x"E1",
     x"E1",
     x"E1",
     x"E1",
     x"E0",
     x"E0",
     x"E0",
     x"E0",
     x"DF",
     x"DF",
     x"DF",
     x"DF",
     x"DE",
     x"DE",
     x"DE",
     x"DE",
     x"DD",
     x"DD",
     x"DD",
     x"DD",
     x"DC",
     x"DC",
     x"DC",
     x"DC",
     x"DB",
     x"DB",
     x"DB",
     x"DB",
     x"DA",
     x"DA",
     x"DA",
     x"DA",
     x"D9",
     x"D9",
     x"D9",
     x"D9",
     x"D8",
     x"D8",
     x"D8",
     x"D7",
     x"D7",
     x"D7",
     x"D7",
     x"D6",
     x"D6",
     x"D6",
     x"D6",
     x"D5",
     x"D5",
     x"D5",
     x"D5",
     x"D4",
     x"D4",
     x"D4",
     x"D3",
     x"D3",
     x"D3",
     x"D3",
     x"D2",
     x"D2",
     x"D2",
     x"D1",
     x"D1",
     x"D1",
     x"D1",
     x"D0",
     x"D0",
     x"D0",
     x"CF",
     x"CF",
     x"CF",
     x"CF",
     x"CE",
     x"CE",
     x"CE",
     x"CD",
     x"CD",
     x"CD",
     x"CC",
     x"CC",
     x"CC",
     x"CC",
     x"CB",
     x"CB",
     x"CB",
     x"CA",
     x"CA",
     x"CA",
     x"C9",
     x"C9",
     x"C9",
     x"C9",
     x"C8",
     x"C8",
     x"C8",
     x"C7",
     x"C7",
     x"C7",
     x"C6",
     x"C6",
     x"C6",
     x"C5",
     x"C5",
     x"C5",
     x"C5",
     x"C4",
     x"C4",
     x"C4",
     x"C3",
     x"C3",
     x"C3",
     x"C2",
     x"C2",
     x"C2",
     x"C1",
     x"C1",
     x"C1",
     x"C0",
     x"C0",
     x"C0",
     x"BF",
     x"BF",
     x"BF",
     x"BE",
     x"BE",
     x"BE",
     x"BD",
     x"BD",
     x"BD",
     x"BC",
     x"BC",
     x"BC",
     x"BB",
     x"BB",
     x"BB",
     x"BA",
     x"BA",
     x"BA",
     x"B9",
     x"B9",
     x"B9",
     x"B8",
     x"B8",
     x"B8",
     x"B7",
     x"B7",
     x"B7",
     x"B6",
     x"B6",
     x"B6",
     x"B5",
     x"B5",
     x"B5",
     x"B4",
     x"B4",
     x"B4",
     x"B3",
     x"B3",
     x"B3",
     x"B2",
     x"B2",
     x"B2",
     x"B1",
     x"B1",
     x"B1",
     x"B0",
     x"B0",
     x"B0",
     x"AF",
     x"AF",
     x"AE",
     x"AE",
     x"AE",
     x"AD",
     x"AD",
     x"AD",
     x"AC",
     x"AC",
     x"AC",
     x"AB",
     x"AB",
     x"AB",
     x"AA",
     x"AA",
     x"A9",
     x"A9",
     x"A9",
     x"A8",
     x"A8",
     x"A8",
     x"A7",
     x"A7",
     x"A7",
     x"A6",
     x"A6",
     x"A6",
     x"A5",
     x"A5",
     x"A4",
     x"A4",
     x"A4",
     x"A3",
     x"A3",
     x"A3",
     x"A2",
     x"A2",
     x"A2",
     x"A1",
     x"A1",
     x"A0",
     x"A0",
     x"A0",
     x"9F",
     x"9F",
     x"9F",
     x"9E",
     x"9E",
     x"9D",
     x"9D",
     x"9D",
     x"9C",
     x"9C",
     x"9C",
     x"9B",
     x"9B",
     x"9B",
     x"9A",
     x"9A",
     x"99",
     x"99",
     x"99",
     x"98",
     x"98",
     x"98",
     x"97",
     x"97",
     x"96",
     x"96",
     x"96",
     x"95",
     x"95",
     x"95",
     x"94",
     x"94",
     x"93",
     x"93",
     x"93",
     x"92",
     x"92",
     x"92",
     x"91",
     x"91",
     x"90",
     x"90",
     x"90",
     x"8F",
     x"8F",
     x"8F",
     x"8E",
     x"8E",
     x"8D",
     x"8D",
     x"8D",
     x"8C",
     x"8C",
     x"8C",
     x"8B",
     x"8B",
     x"8A",
     x"8A",
     x"8A",
     x"89",
     x"89",
     x"89",
     x"88",
     x"88",
     x"87",
     x"87",
     x"87",
     x"86",
     x"86",
     x"85",
     x"85",
     x"85",
     x"84",
     x"84",
     x"84",
     x"83",
     x"83",
     x"82",
     x"82",
     x"82",
     x"81",
     x"81",
     x"81",
     x"80",
     x"80",
     x"7F",
     x"7F",
     x"7F",
     x"7E",
     x"7E",
     x"7D",
     x"7D",
     x"7D",
     x"7C",
     x"7C",
     x"7C",
     x"7B",
     x"7B",
     x"7A",
     x"7A",
     x"7A",
     x"79",
     x"79",
     x"79",
     x"78",
     x"78",
     x"77",
     x"77",
     x"77",
     x"76",
     x"76",
     x"75",
     x"75",
     x"75",
     x"74",
     x"74",
     x"74",
     x"73",
     x"73",
     x"72",
     x"72",
     x"72",
     x"71",
     x"71",
     x"71",
     x"70",
     x"70",
     x"6F",
     x"6F",
     x"6F",
     x"6E",
     x"6E",
     x"6E",
     x"6D",
     x"6D",
     x"6C",
     x"6C",
     x"6C",
     x"6B",
     x"6B",
     x"6B",
     x"6A",
     x"6A",
     x"69",
     x"69",
     x"69",
     x"68",
     x"68",
     x"68",
     x"67",
     x"67",
     x"66",
     x"66",
     x"66",
     x"65",
     x"65",
     x"65",
     x"64",
     x"64",
     x"63",
     x"63",
     x"63",
     x"62",
     x"62",
     x"62",
     x"61",
     x"61",
     x"61",
     x"60",
     x"60",
     x"5F",
     x"5F",
     x"5F",
     x"5E",
     x"5E",
     x"5E",
     x"5D",
     x"5D",
     x"5C",
     x"5C",
     x"5C",
     x"5B",
     x"5B",
     x"5B",
     x"5A",
     x"5A",
     x"5A",
     x"59",
     x"59",
     x"58",
     x"58",
     x"58",
     x"57",
     x"57",
     x"57",
     x"56",
     x"56",
     x"56",
     x"55",
     x"55",
     x"55",
     x"54",
     x"54",
     x"53",
     x"53",
     x"53",
     x"52",
     x"52",
     x"52",
     x"51",
     x"51",
     x"51",
     x"50",
     x"50",
     x"50",
     x"4F",
     x"4F",
     x"4E",
     x"4E",
     x"4E",
     x"4D",
     x"4D",
     x"4D",
     x"4C",
     x"4C",
     x"4C",
     x"4B",
     x"4B",
     x"4B",
     x"4A",
     x"4A",
     x"4A",
     x"49",
     x"49",
     x"49",
     x"48",
     x"48",
     x"48",
     x"47",
     x"47",
     x"47",
     x"46",
     x"46",
     x"46",
     x"45",
     x"45",
     x"45",
     x"44",
     x"44",
     x"44",
     x"43",
     x"43",
     x"43",
     x"42",
     x"42",
     x"42",
     x"41",
     x"41",
     x"41",
     x"40",
     x"40",
     x"40",
     x"3F",
     x"3F",
     x"3F",
     x"3E",
     x"3E",
     x"3E",
     x"3D",
     x"3D",
     x"3D",
     x"3C",
     x"3C",
     x"3C",
     x"3B",
     x"3B",
     x"3B",
     x"3A",
     x"3A",
     x"3A",
     x"39",
     x"39",
     x"39",
     x"39",
     x"38",
     x"38",
     x"38",
     x"37",
     x"37",
     x"37",
     x"36",
     x"36",
     x"36",
     x"35",
     x"35",
     x"35",
     x"35",
     x"34",
     x"34",
     x"34",
     x"33",
     x"33",
     x"33",
     x"32",
     x"32",
     x"32",
     x"32",
     x"31",
     x"31",
     x"31",
     x"30",
     x"30",
     x"30",
     x"2F",
     x"2F",
     x"2F",
     x"2F",
     x"2E",
     x"2E",
     x"2E",
     x"2D",
     x"2D",
     x"2D",
     x"2D",
     x"2C",
     x"2C",
     x"2C",
     x"2B",
     x"2B",
     x"2B",
     x"2B",
     x"2A",
     x"2A",
     x"2A",
     x"29",
     x"29",
     x"29",
     x"29",
     x"28",
     x"28",
     x"28",
     x"28",
     x"27",
     x"27",
     x"27",
     x"27",
     x"26",
     x"26",
     x"26",
     x"25",
     x"25",
     x"25",
     x"25",
     x"24",
     x"24",
     x"24",
     x"24",
     x"23",
     x"23",
     x"23",
     x"23",
     x"22",
     x"22",
     x"22",
     x"22",
     x"21",
     x"21",
     x"21",
     x"21",
     x"20",
     x"20",
     x"20",
     x"20",
     x"1F",
     x"1F",
     x"1F",
     x"1F",
     x"1E",
     x"1E",
     x"1E",
     x"1E",
     x"1D",
     x"1D",
     x"1D",
     x"1D",
     x"1D",
     x"1C",
     x"1C",
     x"1C",
     x"1C",
     x"1B",
     x"1B",
     x"1B",
     x"1B",
     x"1B",
     x"1A",
     x"1A",
     x"1A",
     x"1A",
     x"19",
     x"19",
     x"19",
     x"19",
     x"19",
     x"18",
     x"18",
     x"18",
     x"18",
     x"17",
     x"17",
     x"17",
     x"17",
     x"17",
     x"16",
     x"16",
     x"16",
     x"16",
     x"16",
     x"15",
     x"15",
     x"15",
     x"15",
     x"15",
     x"14",
     x"14",
     x"14",
     x"14",
     x"14",
     x"13",
     x"13",
     x"13",
     x"13",
     x"13",
     x"13",
     x"12",
     x"12",
     x"12",
     x"12",
     x"12",
     x"11",
     x"11",
     x"11",
     x"11",
     x"11",
     x"11",
     x"10",
     x"10",
     x"10",
     x"10",
     x"10",
     x"10",
     x"0F",
     x"0F",
     x"0F",
     x"0F",
     x"0F",
     x"0F",
     x"0E",
     x"0E",
     x"0E",
     x"0E",
     x"0E",
     x"0E",
     x"0D",
     x"0D",
     x"0D",
     x"0D",
     x"0D",
     x"0D",
     x"0D",
     x"0C",
     x"0C",
     x"0C",
     x"0C",
     x"0C",
     x"0C",
     x"0C",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0A",
     x"0A",
     x"0A",
     x"0A",
     x"0A",
     x"0A",
     x"0A",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"03",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"04",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"05",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"06",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"07",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"08",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"09",
     x"0A",
     x"0A",
     x"0A",
     x"0A",
     x"0A",
     x"0A",
     x"0A",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0B",
     x"0C",
     x"0C",
     x"0C",
     x"0C",
     x"0C",
     x"0C",
     x"0C",
     x"0D",
     x"0D",
     x"0D",
     x"0D",
     x"0D",
     x"0D",
     x"0D",
     x"0E",
     x"0E",
     x"0E",
     x"0E",
     x"0E",
     x"0E",
     x"0F",
     x"0F",
     x"0F",
     x"0F",
     x"0F",
     x"0F",
     x"10",
     x"10",
     x"10",
     x"10",
     x"10",
     x"10",
     x"11",
     x"11",
     x"11",
     x"11",
     x"11",
     x"11",
     x"12",
     x"12",
     x"12",
     x"12",
     x"12",
     x"13",
     x"13",
     x"13",
     x"13",
     x"13",
     x"13",
     x"14",
     x"14",
     x"14",
     x"14",
     x"14",
     x"15",
     x"15",
     x"15",
     x"15",
     x"15",
     x"16",
     x"16",
     x"16",
     x"16",
     x"16",
     x"17",
     x"17",
     x"17",
     x"17",
     x"17",
     x"18",
     x"18",
     x"18",
     x"18",
     x"19",
     x"19",
     x"19",
     x"19",
     x"19",
     x"1A",
     x"1A",
     x"1A",
     x"1A",
     x"1B",
     x"1B",
     x"1B",
     x"1B",
     x"1B",
     x"1C",
     x"1C",
     x"1C",
     x"1C",
     x"1D",
     x"1D",
     x"1D",
     x"1D",
     x"1D",
     x"1E",
     x"1E",
     x"1E",
     x"1E",
     x"1F",
     x"1F",
     x"1F",
     x"1F",
     x"20",
     x"20",
     x"20",
     x"20",
     x"21",
     x"21",
     x"21",
     x"21",
     x"22",
     x"22",
     x"22",
     x"22",
     x"23",
     x"23",
     x"23",
     x"23",
     x"24",
     x"24",
     x"24",
     x"24",
     x"25",
     x"25",
     x"25",
     x"25",
     x"26",
     x"26",
     x"26",
     x"27",
     x"27",
     x"27",
     x"27",
     x"28",
     x"28",
     x"28",
     x"28",
     x"29",
     x"29",
     x"29",
     x"29",
     x"2A",
     x"2A",
     x"2A",
     x"2B",
     x"2B",
     x"2B",
     x"2B",
     x"2C",
     x"2C",
     x"2C",
     x"2D",
     x"2D",
     x"2D",
     x"2D",
     x"2E",
     x"2E",
     x"2E",
     x"2F",
     x"2F",
     x"2F",
     x"2F",
     x"30",
     x"30",
     x"30",
     x"31",
     x"31",
     x"31",
     x"32",
     x"32",
     x"32",
     x"32",
     x"33",
     x"33",
     x"33",
     x"34",
     x"34",
     x"34",
     x"35",
     x"35",
     x"35",
     x"35",
     x"36",
     x"36",
     x"36",
     x"37",
     x"37",
     x"37",
     x"38",
     x"38",
     x"38",
     x"39",
     x"39",
     x"39",
     x"39",
     x"3A",
     x"3A",
     x"3A",
     x"3B",
     x"3B",
     x"3B",
     x"3C",
     x"3C",
     x"3C",
     x"3D",
     x"3D",
     x"3D",
     x"3E",
     x"3E",
     x"3E",
     x"3F",
     x"3F",
     x"3F",
     x"40",
     x"40",
     x"40",
     x"41",
     x"41",
     x"41",
     x"42",
     x"42",
     x"42",
     x"43",
     x"43",
     x"43",
     x"44",
     x"44",
     x"44",
     x"45",
     x"45",
     x"45",
     x"46",
     x"46",
     x"46",
     x"47",
     x"47",
     x"47",
     x"48",
     x"48",
     x"48",
     x"49",
     x"49",
     x"49",
     x"4A",
     x"4A",
     x"4A",
     x"4B",
     x"4B",
     x"4B",
     x"4C",
     x"4C",
     x"4C",
     x"4D",
     x"4D",
     x"4D",
     x"4E",
     x"4E",
     x"4E",
     x"4F",
     x"4F",
     x"50",
     x"50",
     x"50",
     x"51",
     x"51",
     x"51",
     x"52",
     x"52",
     x"52",
     x"53",
     x"53",
     x"53",
     x"54",
     x"54",
     x"55",
     x"55",
     x"55",
     x"56",
     x"56",
     x"56",
     x"57",
     x"57",
     x"57",
     x"58",
     x"58",
     x"58",
     x"59",
     x"59",
     x"5A",
     x"5A",
     x"5A",
     x"5B",
     x"5B",
     x"5B",
     x"5C",
     x"5C",
     x"5C",
     x"5D",
     x"5D",
     x"5E",
     x"5E",
     x"5E",
     x"5F",
     x"5F",
     x"5F",
     x"60",
     x"60",
     x"61",
     x"61",
     x"61",
     x"62",
     x"62",
     x"62",
     x"63",
     x"63",
     x"63",
     x"64",
     x"64",
     x"65",
     x"65",
     x"65",
     x"66",
     x"66",
     x"66",
     x"67",
     x"67",
     x"68",
     x"68",
     x"68",
     x"69",
     x"69",
     x"69",
     x"6A",
     x"6A",
     x"6B",
     x"6B",
     x"6B",
     x"6C",
     x"6C",
     x"6C",
     x"6D",
     x"6D",
     x"6E",
     x"6E",
     x"6E",
     x"6F",
     x"6F",
     x"6F",
     x"70",
     x"70",
     x"71",
     x"71",
     x"71",
     x"72",
     x"72",
     x"72",
     x"73",
     x"73",
     x"74",
     x"74",
     x"74",
     x"75",
     x"75",
     x"75",
     x"76",
     x"76",
     x"77",
     x"77",
     x"77",
     x"78",
     x"78",
     x"79",
     x"79",
     x"79",
     x"7A",
     x"7A",
     x"7A",
     x"7B",
     x"7B",
     x"7C",
     x"7C",
     x"7C",
     x"7D",
     x"7D",
     x"7D",
     x"7E",
     x"7F"
    );
    signal data_counter : std_logic_vector(11 downto 0):=(others => '0');
    signal data_d       : std_logic_vector(7 downto 0);

begin

addr_proc :
  process(clk)
  begin
    if rising_edge(clk) then
      if rst = '1' then
        data_counter <= (others => '0');
      else
        if ((start = '1') and (data_counter = 0)) then 
          data_counter <= data_counter + 1;
        end if;
        if ((data_counter > 0) and (data_counter(data_counter'length - 1) = '0')) then
          data_counter <= data_counter + 1;
        end if;
      end if;
      data <= sin_form(to_integer(unsigned(data_counter(data_counter'length - 2 downto 0))));
      addr <= data_counter(addr'length - 1 downto 0);
      wr_en <= not(data_counter(data_counter'length - 1));
    end if;
  end process;



end Behavioral;
